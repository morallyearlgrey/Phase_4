module INSTRUCTION_MEMORY (
    input iRdAddr,
    output [31:0] oInstr
);
    
endmodule