module DATA_MEMORY (
    input [31:0] iAddress,
    input [31:0] iWriteData,
    input [2:0] iFunct3,
    input iMemWrite,
    input iMemRead,
    output reg [31:0] oReadData
);
    
endmodule