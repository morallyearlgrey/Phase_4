module BRANCH_JUMP (
    input iBranch,
    input iJump,
    input iZero,
    input [31:0] iOffset,
    input [31:0] iPc,
    input [31:0] iRs1,
    input iPcSrc,
    output [31:0] oPc
);
    
endmodule